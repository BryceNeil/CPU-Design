module or_new (input x, y, output z);

assign z = x | y;

	endmodule