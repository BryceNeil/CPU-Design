`timescale 1ns/1ps

module register_tb;

//module register (BusMuxOut, clr, clk, Rin, BusMuxIn_R);

reg reg_in, clk ;

endmodule